module orGate
#(parameter N=4)

(input logic [N-1:0] a,
 input logic [N-1:0] b,
 output logic [N-1:0] result);
 

    always_comb begin
        result = a | b;
    end

endmodule
