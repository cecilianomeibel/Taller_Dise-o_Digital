module moduleN
#(parameter N=4)

( input logic [N-1:0] dividend,  //dividendo
  input logic [N-1:0] divider,   //divisor
  output logic [N-1:0] remainder //resto
);


always_comb begin

remainder = dividend % divider;

end
endmodule
