module dividerN

#(parameter N = 4) 

( input logic [N-1:0] dividend, //dividendo
  input logic [N-1:0] divider, // divisor
  output logic [N-1:0] quotient //cociente
);

always_comb begin

quotient= dividend/divider;

end 

endmodule